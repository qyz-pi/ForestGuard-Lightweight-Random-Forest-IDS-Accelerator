`ifndef RF_ADDRS_VH
`define RF_ADDRS_VH

`define RF_NUM_TREES 6
`define RF_NODE_WIDTH 36

localparam integer BASE0 = 0;
localparam integer BASE1 = 311;
localparam integer BASE2 = 680;
localparam integer BASE3 = 985;
localparam integer BASE4 = 1332;
localparam integer BASE5 = 1635;

`endif // RF_ADDRS_VH
